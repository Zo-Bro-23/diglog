module morse(inout [33:0] GPIO, input CLOCK_50, output [17:0] LEDR);
	assign LEDR = GPIO[25:17];
	assign GPIO[33:26] = GPIO[25:18];
	interpret(CLOCK_50, GPIO[25:18], GPIO[17], GPIO[2:0], GPIO[6:4], GPIO[11:8], GPIO[12], GPIO[13], GPIO[14], GPIO[3], GPIO[15], GPIO[7]);
endmodule

module interpret(input CLOCK, input [7:0] letter, input ardCLK, output reg [2:0] RGB1, output reg [2:0] RGB2, output reg [3:0] addr, output reg CLK, LAT, OE, output GND1, GND2, GND3);
	assign GND1 = 0;
	assign GND2 = 0;
	assign GND3 = 0;
		
	reg clk;
	
	reg [24:0] clkcounter = 0;
	reg [24:0] rowcounter = 8025;
	reg [24:0] addrcounter = 0;

	reg [223:0] store1 = 224'b00000000011111100100001001000010010000100100001001000010011111100011110000111110001111000011111000111100010000100100001000000010010000100111100000111100010000100011110001111110011111100001111000111100001111100001100000000000;
	reg [223:0] store2 = 224'b00000000010000000100001001000010010000100100001001000010000010000100001001000010010000100100001001000010010001100110011000000010001000100010000000001000010000100100001000000010000000100010001001000010010000100010010000000000;
	reg [223:0] store3 = 224'b00000000001000000010010000100100010000100100001001000010000010000000001001000010010000100100001001000010010010100101101000000010000100100010000000001000010000100000001000000010000000100100001000000010010000100100001000000000;
	reg [223:0] store4 = 224'b00000000000100000001100000011000010000100100001001000010000010000011110000111110010000100011111001000010010100100101101000000010000011100010000000001000011111100000001000111110001111100100001000000010001111100100001000000000;
	reg [223:0] store5 = 224'b00000000000010000000100000011000010110100100001001000010000010000100000000010010010000100000001001000010011000100100001000000010000100100010000000001000010000100111001000000010000000100100001000000010010000100111111000000000;
	reg [223:0] store6 = 224'b00001110000001000000100000100100010110100100001001000010000010000100000000100010010100100000001001000010010000100100001000000010001000100010001000001000010000100100001000000010000000100100001000000010010000100100001000000000;
	reg [223:0] store7 = 224'b00001110000000100000100001000010011001100010010001000010000010000100001001000010001000100000001001000010010000100100001000000010010000100010001000001000010000100100001000000010000000100010001001000010010000100100001000000000;
	reg [223:0] store8 = 224'b00001110011111100000100001000010010000100001100000111100000010000011110001000010010111000000001000111100010000100100001001111110010000100001110000111100010000100011110000000010011111100001111000111100001111100100001000000000;
	
	reg [63:0] symb1 = 64'b0001100000000000000000000000000000001111111100000000000000000000;
	reg [63:0] symb2 = 64'b0011100000000000000000000000000000001111111100000000000000000000;
	reg [63:0] symb3 = 64'b0111100000000000000000000000000000001111111100000000000000000000;
	reg [63:0] symb4 = 64'b1111111111111111111111111111111100001111111100000000000000000000;
	reg [63:0] symb5 = 64'b1111111111111111111111111111111100001111111100000000000000000000;
	reg [63:0] symb6 = 64'b0111100000000000000000000000000000001111111100000000000000000000;
	reg [63:0] symb7 = 64'b0011100000000000000000000000000000001111111100000000000000000000;
	reg [63:0] symb8 = 64'b0001100000000000000000000000000000001111111100000000000000000000;
	
	reg [1791:0] store;
	reg [511:0] symb;
	
	reg [511:0] row1;
	reg [511:0] row2;
	
	reg [5:0] i;
		
	always @ (*) begin
		store <= {store8, store7, store6, store5, store4, store3, store2, store1};
		symb <= {symb8, symb7, symb6, symb5, symb4, symb3, symb2, symb1};
	end
	
	always @ (posedge CLOCK) begin
		clkcounter = clkcounter + 1;
		if (clkcounter == 1) begin
			clkcounter = 0;
			clk = !clk;
			if (rowcounter <= 63) CLK = clk;
			else CLK = 0;
		end
	end
	
	always @ (posedge clk) begin
		if (rowcounter <= 63) begin
			if (addrcounter <= 11 && addrcounter >= 4) begin
				RGB1 <= {3{row1[(addrcounter - 4) * 64 + rowcounter]}};
				RGB2 <= {3{row2[(addrcounter - 4) * 64 + rowcounter]}};
			end
			else begin
				RGB1 <= 3'b000;
				RGB2 <= 3'b000;
			end
		end
		if (rowcounter == 500) OE <= 0;
		if (rowcounter == 550) LAT <= 1;
		if (rowcounter == 600) LAT <= 0;
		if (rowcounter == 650) OE <= 1;
		rowcounter <= rowcounter + 1;
		if (rowcounter == 8000) begin
			addr <= addr + 1;
			addrcounter[3:0] <= addr + 2;
		end
		if (rowcounter == 8050) rowcounter <= 0;
end
			
	always @ (posedge ardCLK) begin
		for (i = 0; i < 8; i = i + 1) begin
			if(letter >= 29) begin
				row1[(i * 64) +: 64] <= {{24{1'b0}}, symb[(i * 64) + ((letter - 29) * 16) +: 16], {24{1'b0}}};
				row2 <= {64{3'b000}};
			end
			else begin
				row2[(i * 64) +: 56] <= row2[(i * 64 + 8) +: 56];
				row2[(i * 64 + 56) +: 8] <= {store[(i * 224) + ((letter - 1) * 8) +: 8]}; // Index of 0 does not work with Arduino
				row1 <= {64{3'b000}};
			end
		end
	end
endmodule
